// QSYS_CORE_tb.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module QSYS_CORE_tb (
	);

	wire          qsys_core_inst_clk_bfm_clk_clk;                    // QSYS_CORE_inst_clk_bfm:clk -> [QSYS_CORE_inst:clk_clk, QSYS_CORE_inst_reset_bfm:clk]
	wire    [1:0] qsys_core_inst_axi4_mst_128_bfm_conduit_awburst;   // QSYS_CORE_inst_axi4_mst_128_bfm:sig_awburst -> QSYS_CORE_inst:axi4_mst_128_awburst
	wire   [31:0] qsys_core_inst_axi4_mst_128_bfm_conduit_awaddr;    // QSYS_CORE_inst_axi4_mst_128_bfm:sig_awaddr -> QSYS_CORE_inst:axi4_mst_128_awaddr
	wire    [7:0] qsys_core_inst_axi4_mst_128_bfm_conduit_arlen;     // QSYS_CORE_inst_axi4_mst_128_bfm:sig_arlen -> QSYS_CORE_inst:axi4_mst_128_arlen
	wire          qsys_core_inst_axi4_mst_128_arready;               // QSYS_CORE_inst:axi4_mst_128_arready -> QSYS_CORE_inst_axi4_mst_128_bfm:sig_arready
	wire  [127:0] qsys_core_inst_axi4_mst_128_rdata;                 // QSYS_CORE_inst:axi4_mst_128_rdata -> QSYS_CORE_inst_axi4_mst_128_bfm:sig_rdata
	wire          qsys_core_inst_axi4_mst_128_wready;                // QSYS_CORE_inst:axi4_mst_128_wready -> QSYS_CORE_inst_axi4_mst_128_bfm:sig_wready
	wire    [1:0] qsys_core_inst_axi4_mst_128_bfm_conduit_arburst;   // QSYS_CORE_inst_axi4_mst_128_bfm:sig_arburst -> QSYS_CORE_inst:axi4_mst_128_arburst
	wire          qsys_core_inst_axi4_mst_128_awready;               // QSYS_CORE_inst:axi4_mst_128_awready -> QSYS_CORE_inst_axi4_mst_128_bfm:sig_awready
	wire    [0:0] qsys_core_inst_axi4_mst_128_bfm_conduit_rready;    // QSYS_CORE_inst_axi4_mst_128_bfm:sig_rready -> QSYS_CORE_inst:axi4_mst_128_rready
	wire    [2:0] qsys_core_inst_axi4_mst_128_bfm_conduit_arsize;    // QSYS_CORE_inst_axi4_mst_128_bfm:sig_arsize -> QSYS_CORE_inst:axi4_mst_128_arsize
	wire    [7:0] qsys_core_inst_axi4_mst_128_bfm_conduit_awlen;     // QSYS_CORE_inst_axi4_mst_128_bfm:sig_awlen -> QSYS_CORE_inst:axi4_mst_128_awlen
	wire    [0:0] qsys_core_inst_axi4_mst_128_bfm_conduit_bready;    // QSYS_CORE_inst_axi4_mst_128_bfm:sig_bready -> QSYS_CORE_inst:axi4_mst_128_bready
	wire          qsys_core_inst_axi4_mst_128_rlast;                 // QSYS_CORE_inst:axi4_mst_128_rlast -> QSYS_CORE_inst_axi4_mst_128_bfm:sig_rlast
	wire    [0:0] qsys_core_inst_axi4_mst_128_bfm_conduit_wlast;     // QSYS_CORE_inst_axi4_mst_128_bfm:sig_wlast -> QSYS_CORE_inst:axi4_mst_128_wlast
	wire   [31:0] qsys_core_inst_axi4_mst_128_bfm_conduit_araddr;    // QSYS_CORE_inst_axi4_mst_128_bfm:sig_araddr -> QSYS_CORE_inst:axi4_mst_128_araddr
	wire    [0:0] qsys_core_inst_axi4_mst_128_bfm_conduit_wvalid;    // QSYS_CORE_inst_axi4_mst_128_bfm:sig_wvalid -> QSYS_CORE_inst:axi4_mst_128_wvalid
	wire    [2:0] qsys_core_inst_axi4_mst_128_bfm_conduit_arprot;    // QSYS_CORE_inst_axi4_mst_128_bfm:sig_arprot -> QSYS_CORE_inst:axi4_mst_128_arprot
	wire    [0:0] qsys_core_inst_axi4_mst_128_bfm_conduit_arvalid;   // QSYS_CORE_inst_axi4_mst_128_bfm:sig_arvalid -> QSYS_CORE_inst:axi4_mst_128_arvalid
	wire    [2:0] qsys_core_inst_axi4_mst_128_bfm_conduit_awprot;    // QSYS_CORE_inst_axi4_mst_128_bfm:sig_awprot -> QSYS_CORE_inst:axi4_mst_128_awprot
	wire  [127:0] qsys_core_inst_axi4_mst_128_bfm_conduit_wdata;     // QSYS_CORE_inst_axi4_mst_128_bfm:sig_wdata -> QSYS_CORE_inst:axi4_mst_128_wdata
	wire          qsys_core_inst_axi4_mst_128_bvalid;                // QSYS_CORE_inst:axi4_mst_128_bvalid -> QSYS_CORE_inst_axi4_mst_128_bfm:sig_bvalid
	wire    [2:0] qsys_core_inst_axi4_mst_128_bfm_conduit_awsize;    // QSYS_CORE_inst_axi4_mst_128_bfm:sig_awsize -> QSYS_CORE_inst:axi4_mst_128_awsize
	wire    [0:0] qsys_core_inst_axi4_mst_128_bfm_conduit_awvalid;   // QSYS_CORE_inst_axi4_mst_128_bfm:sig_awvalid -> QSYS_CORE_inst:axi4_mst_128_awvalid
	wire          qsys_core_inst_axi4_mst_128_rvalid;                // QSYS_CORE_inst:axi4_mst_128_rvalid -> QSYS_CORE_inst_axi4_mst_128_bfm:sig_rvalid
	wire          qsys_core_inst_axi4_mst_128_reset_reset;           // QSYS_CORE_inst:axi4_mst_128_reset_reset -> QSYS_CORE_inst_axi4_mst_128_reset_bfm:sig_reset
	wire    [1:0] qsys_core_inst_axi4_mst_16_bfm_conduit_awburst;    // QSYS_CORE_inst_axi4_mst_16_bfm:sig_awburst -> QSYS_CORE_inst:axi4_mst_16_awburst
	wire   [31:0] qsys_core_inst_axi4_mst_16_bfm_conduit_awaddr;     // QSYS_CORE_inst_axi4_mst_16_bfm:sig_awaddr -> QSYS_CORE_inst:axi4_mst_16_awaddr
	wire    [7:0] qsys_core_inst_axi4_mst_16_bfm_conduit_arlen;      // QSYS_CORE_inst_axi4_mst_16_bfm:sig_arlen -> QSYS_CORE_inst:axi4_mst_16_arlen
	wire          qsys_core_inst_axi4_mst_16_arready;                // QSYS_CORE_inst:axi4_mst_16_arready -> QSYS_CORE_inst_axi4_mst_16_bfm:sig_arready
	wire   [15:0] qsys_core_inst_axi4_mst_16_rdata;                  // QSYS_CORE_inst:axi4_mst_16_rdata -> QSYS_CORE_inst_axi4_mst_16_bfm:sig_rdata
	wire          qsys_core_inst_axi4_mst_16_wready;                 // QSYS_CORE_inst:axi4_mst_16_wready -> QSYS_CORE_inst_axi4_mst_16_bfm:sig_wready
	wire    [1:0] qsys_core_inst_axi4_mst_16_bfm_conduit_arburst;    // QSYS_CORE_inst_axi4_mst_16_bfm:sig_arburst -> QSYS_CORE_inst:axi4_mst_16_arburst
	wire          qsys_core_inst_axi4_mst_16_awready;                // QSYS_CORE_inst:axi4_mst_16_awready -> QSYS_CORE_inst_axi4_mst_16_bfm:sig_awready
	wire    [0:0] qsys_core_inst_axi4_mst_16_bfm_conduit_rready;     // QSYS_CORE_inst_axi4_mst_16_bfm:sig_rready -> QSYS_CORE_inst:axi4_mst_16_rready
	wire    [2:0] qsys_core_inst_axi4_mst_16_bfm_conduit_arsize;     // QSYS_CORE_inst_axi4_mst_16_bfm:sig_arsize -> QSYS_CORE_inst:axi4_mst_16_arsize
	wire    [7:0] qsys_core_inst_axi4_mst_16_bfm_conduit_awlen;      // QSYS_CORE_inst_axi4_mst_16_bfm:sig_awlen -> QSYS_CORE_inst:axi4_mst_16_awlen
	wire    [0:0] qsys_core_inst_axi4_mst_16_bfm_conduit_bready;     // QSYS_CORE_inst_axi4_mst_16_bfm:sig_bready -> QSYS_CORE_inst:axi4_mst_16_bready
	wire          qsys_core_inst_axi4_mst_16_rlast;                  // QSYS_CORE_inst:axi4_mst_16_rlast -> QSYS_CORE_inst_axi4_mst_16_bfm:sig_rlast
	wire    [0:0] qsys_core_inst_axi4_mst_16_bfm_conduit_wlast;      // QSYS_CORE_inst_axi4_mst_16_bfm:sig_wlast -> QSYS_CORE_inst:axi4_mst_16_wlast
	wire   [31:0] qsys_core_inst_axi4_mst_16_bfm_conduit_araddr;     // QSYS_CORE_inst_axi4_mst_16_bfm:sig_araddr -> QSYS_CORE_inst:axi4_mst_16_araddr
	wire    [0:0] qsys_core_inst_axi4_mst_16_bfm_conduit_wvalid;     // QSYS_CORE_inst_axi4_mst_16_bfm:sig_wvalid -> QSYS_CORE_inst:axi4_mst_16_wvalid
	wire    [2:0] qsys_core_inst_axi4_mst_16_bfm_conduit_arprot;     // QSYS_CORE_inst_axi4_mst_16_bfm:sig_arprot -> QSYS_CORE_inst:axi4_mst_16_arprot
	wire    [0:0] qsys_core_inst_axi4_mst_16_bfm_conduit_arvalid;    // QSYS_CORE_inst_axi4_mst_16_bfm:sig_arvalid -> QSYS_CORE_inst:axi4_mst_16_arvalid
	wire    [2:0] qsys_core_inst_axi4_mst_16_bfm_conduit_awprot;     // QSYS_CORE_inst_axi4_mst_16_bfm:sig_awprot -> QSYS_CORE_inst:axi4_mst_16_awprot
	wire   [15:0] qsys_core_inst_axi4_mst_16_bfm_conduit_wdata;      // QSYS_CORE_inst_axi4_mst_16_bfm:sig_wdata -> QSYS_CORE_inst:axi4_mst_16_wdata
	wire          qsys_core_inst_axi4_mst_16_bvalid;                 // QSYS_CORE_inst:axi4_mst_16_bvalid -> QSYS_CORE_inst_axi4_mst_16_bfm:sig_bvalid
	wire    [2:0] qsys_core_inst_axi4_mst_16_bfm_conduit_awsize;     // QSYS_CORE_inst_axi4_mst_16_bfm:sig_awsize -> QSYS_CORE_inst:axi4_mst_16_awsize
	wire    [0:0] qsys_core_inst_axi4_mst_16_bfm_conduit_awvalid;    // QSYS_CORE_inst_axi4_mst_16_bfm:sig_awvalid -> QSYS_CORE_inst:axi4_mst_16_awvalid
	wire          qsys_core_inst_axi4_mst_16_rvalid;                 // QSYS_CORE_inst:axi4_mst_16_rvalid -> QSYS_CORE_inst_axi4_mst_16_bfm:sig_rvalid
	wire          qsys_core_inst_axi4_mst_16_reset_reset;            // QSYS_CORE_inst:axi4_mst_16_reset_reset -> QSYS_CORE_inst_axi4_mst_16_reset_bfm:sig_reset
	wire   [15:0] qsys_core_inst_axi4lite_slv_0_awaddr;              // QSYS_CORE_inst:axi4lite_slv_0_awaddr -> QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_awaddr
	wire    [0:0] qsys_core_inst_axi4lite_slv_0_bfm_conduit_arready; // QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_arready -> QSYS_CORE_inst:axi4lite_slv_0_arready
	wire    [1:0] qsys_core_inst_axi4lite_slv_0_bfm_conduit_bresp;   // QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_bresp -> QSYS_CORE_inst:axi4lite_slv_0_bresp
	wire   [31:0] qsys_core_inst_axi4lite_slv_0_bfm_conduit_rdata;   // QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_rdata -> QSYS_CORE_inst:axi4lite_slv_0_rdata
	wire    [0:0] qsys_core_inst_axi4lite_slv_0_bfm_conduit_wready;  // QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_wready -> QSYS_CORE_inst:axi4lite_slv_0_wready
	wire    [3:0] qsys_core_inst_axi4lite_slv_0_wstrb;               // QSYS_CORE_inst:axi4lite_slv_0_wstrb -> QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_wstrb
	wire    [0:0] qsys_core_inst_axi4lite_slv_0_bfm_conduit_awready; // QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_awready -> QSYS_CORE_inst:axi4lite_slv_0_awready
	wire          qsys_core_inst_axi4lite_slv_0_rready;              // QSYS_CORE_inst:axi4lite_slv_0_rready -> QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_rready
	wire          qsys_core_inst_axi4lite_slv_0_bready;              // QSYS_CORE_inst:axi4lite_slv_0_bready -> QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_bready
	wire   [15:0] qsys_core_inst_axi4lite_slv_0_araddr;              // QSYS_CORE_inst:axi4lite_slv_0_araddr -> QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_araddr
	wire          qsys_core_inst_axi4lite_slv_0_wvalid;              // QSYS_CORE_inst:axi4lite_slv_0_wvalid -> QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_wvalid
	wire    [2:0] qsys_core_inst_axi4lite_slv_0_arprot;              // QSYS_CORE_inst:axi4lite_slv_0_arprot -> QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_arprot
	wire    [1:0] qsys_core_inst_axi4lite_slv_0_bfm_conduit_rresp;   // QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_rresp -> QSYS_CORE_inst:axi4lite_slv_0_rresp
	wire          qsys_core_inst_axi4lite_slv_0_arvalid;             // QSYS_CORE_inst:axi4lite_slv_0_arvalid -> QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_arvalid
	wire    [2:0] qsys_core_inst_axi4lite_slv_0_awprot;              // QSYS_CORE_inst:axi4lite_slv_0_awprot -> QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_awprot
	wire   [31:0] qsys_core_inst_axi4lite_slv_0_wdata;               // QSYS_CORE_inst:axi4lite_slv_0_wdata -> QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_wdata
	wire    [0:0] qsys_core_inst_axi4lite_slv_0_bfm_conduit_bvalid;  // QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_bvalid -> QSYS_CORE_inst:axi4lite_slv_0_bvalid
	wire          qsys_core_inst_axi4lite_slv_0_awvalid;             // QSYS_CORE_inst:axi4lite_slv_0_awvalid -> QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_awvalid
	wire    [0:0] qsys_core_inst_axi4lite_slv_0_bfm_conduit_rvalid;  // QSYS_CORE_inst_axi4lite_slv_0_bfm:sig_rvalid -> QSYS_CORE_inst:axi4lite_slv_0_rvalid
	wire          qsys_core_inst_axi4lite_slv_0_reset_reset;         // QSYS_CORE_inst:axi4lite_slv_0_reset_reset -> QSYS_CORE_inst_axi4lite_slv_0_reset_bfm:sig_reset
	wire    [7:0] qsys_core_inst_pio_out_export;                     // QSYS_CORE_inst:pio_out_export -> QSYS_CORE_inst_pio_out_bfm:sig_export
	wire          qsys_core_inst_reset_bfm_reset_reset;              // QSYS_CORE_inst_reset_bfm:reset -> QSYS_CORE_inst:reset_reset_n

	QSYS_CORE qsys_core_inst (
		.axi4_mst_128_awaddr        (32'b0),    //         axi4_mst_128.awaddr
		.axi4_mst_128_awprot        (3'b0),    //                     .awprot
		.axi4_mst_128_awvalid       (1'b0),   //                     .awvalid
		.axi4_mst_128_awready       (),               //                     .awready
		.axi4_mst_128_wdata         (32'b0),     //                     .wdata
		.axi4_mst_128_wlast         (1'b0),     //                     .wlast
		.axi4_mst_128_wvalid        (1'b0),    //                     .wvalid
		.axi4_mst_128_wready        (),                //                     .wready
		.axi4_mst_128_bvalid        (),                //                     .bvalid
		.axi4_mst_128_bready        (1'b0),    //                     .bready
		.axi4_mst_128_araddr        (1'b0),    //                     .araddr
		.axi4_mst_128_arprot        (1'b0),    //                     .arprot
		.axi4_mst_128_arvalid       (1'b0),   //                     .arvalid
		.axi4_mst_128_arready       (),               //                     .arready
		.axi4_mst_128_rdata         (),                 //                     .rdata
		.axi4_mst_128_rvalid        (),                //                     .rvalid
		.axi4_mst_128_rready        (1'b0),    //                     .rready
		.axi4_mst_128_arlen         (1'b0),     //                     .arlen
		.axi4_mst_128_arburst       (1'b0),   //                     .arburst
		.axi4_mst_128_arsize        (1'b0),    //                     .arsize
		.axi4_mst_128_awlen         (1'b0),     //                     .awlen
		.axi4_mst_128_awburst       (1'b0),   //                     .awburst
		.axi4_mst_128_awsize        (1'b0),    //                     .awsize
		.axi4_mst_128_rlast         (),                 //                     .rlast
		.axi4_mst_128_reset_reset   (qsys_core_inst_axi4_mst_128_reset_reset),           //   axi4_mst_128_reset.reset
		.axi4_mst_16_awaddr         (1'b0),     //          axi4_mst_16.awaddr
		.axi4_mst_16_awprot         (1'b0),     //                     .awprot
		.axi4_mst_16_awvalid        (1'b0),    //                     .awvalid
		.axi4_mst_16_awready        (),                //                     .awready
		.axi4_mst_16_wdata          (1'b0),      //                     .wdata
		.axi4_mst_16_wlast          (1'b0),      //                     .wlast
		.axi4_mst_16_wvalid         (1'b0),     //                     .wvalid
		.axi4_mst_16_wready         (),                 //                     .wready
		.axi4_mst_16_bvalid         (),                 //                     .bvalid
		.axi4_mst_16_bready         (1'b0),     //                     .bready
		.axi4_mst_16_araddr         (1'b0),     //                     .araddr
		.axi4_mst_16_arprot         (1'b0),     //                     .arprot
		.axi4_mst_16_arvalid        (1'b0),    //                     .arvalid
		.axi4_mst_16_arready        (),                //                     .arready
		.axi4_mst_16_rdata          (),                  //                     .rdata
		.axi4_mst_16_rvalid         (),                 //                     .rvalid
		.axi4_mst_16_rready         (1'b0),     //                     .rready
		.axi4_mst_16_arlen          (1'b0),      //                     .arlen
		.axi4_mst_16_arburst        (1'b0),    //                     .arburst
		.axi4_mst_16_arsize         (1'b0),     //                     .arsize
		.axi4_mst_16_awlen          (1'b0),      //                     .awlen
		.axi4_mst_16_awburst        (1'b0),    //                     .awburst
		.axi4_mst_16_awsize         (1'b0),     //                     .awsize
		.axi4_mst_16_rlast          (),                  //                     .rlast
		.axi4_mst_16_reset_reset    (qsys_core_inst_axi4_mst_16_reset_reset),            //    axi4_mst_16_reset.reset
		.axi4lite_slv_0_araddr      (),              //       axi4lite_slv_0.araddr
		.axi4lite_slv_0_arready     (1'b0), //                     .arready
		.axi4lite_slv_0_awaddr      (),              //                     .awaddr
		.axi4lite_slv_0_awready     (1'b0), //                     .awready
		.axi4lite_slv_0_arvalid     (),             //                     .arvalid
		.axi4lite_slv_0_awvalid     (),             //                     .awvalid
		.axi4lite_slv_0_rdata       (1'b0),   //                     .rdata
		.axi4lite_slv_0_rready      (),              //                     .rready
		.axi4lite_slv_0_rvalid      (1'b0),  //                     .rvalid
		.axi4lite_slv_0_wdata       (),               //                     .wdata
		.axi4lite_slv_0_wready      (1'b0),  //                     .wready
		.axi4lite_slv_0_wstrb       (),               //                     .wstrb
		.axi4lite_slv_0_wvalid      (),              //                     .wvalid
		.axi4lite_slv_0_arprot      (),              //                     .arprot
		.axi4lite_slv_0_awprot      (),              //                     .awprot
		.axi4lite_slv_0_bready      (),              //                     .bready
		.axi4lite_slv_0_bresp       (1'b0),   //                     .bresp
		.axi4lite_slv_0_bvalid      (1'b0),  //                     .bvalid
		.axi4lite_slv_0_rresp       (1'b0),   //                     .rresp
		.axi4lite_slv_0_reset_reset (),         // axi4lite_slv_0_reset.reset
		.clk_clk                    (qsys_core_inst_clk_bfm_clk_clk),                    //                  clk.clk
		.pio_out_export             (qsys_core_inst_pio_out_export),                     //              pio_out.export
		.reset_reset_n              (qsys_core_inst_reset_bfm_reset_reset)               //                reset.reset_n
	);


    block_t 
//    #(.IDWIDTH(IDWIDTH),
//      .IDNUM  (IDNUM0),
//      .BSIZE  (BSIZE),
//      .DWB    (DWB),
//      .DW     (DW)
//     ) block_t_inst
	block_t block_t_inst (
      .i_clk(qsys_core_inst_clk_bfm_clk_clk),
      .i_rst_n(qsys_core_inst_reset_bfm_reset_reset),
      .rggen_axi4lite_if.slave axi4lite_if(),
      .o_register_0_bit_field_0(),
      .o_register_0_bit_field_1(),
      .o_register_0_bit_field_2(),
      .o_register_1_bit_field_0(),
      .o_register_1_bit_field_1(),
      .o_register_2_bit_field_0(),
      .o_register_3_bit_field_0(),
      .o_register_4_bit_field_0(),
      .o_register_5_bit_field_0(),
      .o_register_6_bit_field_0(),
      .o_register_7_bit_field_0()
	 );

module block_t
  import rggen_rtl_pkg::*;
#(
  parameter int ADDRESS_WIDTH = 5,
  parameter bit PRE_DECODE = 0,
  parameter bit [ADDRESS_WIDTH-1:0] BASE_ADDRESS = '0,
  parameter bit ERROR_STATUS = 0,
  parameter bit [31:0] DEFAULT_READ_DATA = '0,
  parameter int ID_WIDTH = 0,
  parameter bit WRITE_FIRST = 1
)(
  input logic i_clk,
  input logic i_rst_n,
  rggen_axi4lite_if.slave axi4lite_if,
  output logic [3:0] o_register_0_bit_field_0,
  output logic [3:0] o_register_0_bit_field_1,
  output logic o_register_0_bit_field_2,
  output logic [15:0] o_register_1_bit_field_0,
  output logic [15:0] o_register_1_bit_field_1,
  output logic [31:0] o_register_2_bit_field_0,
  output logic [31:0] o_register_3_bit_field_0,
  output logic [31:0] o_register_4_bit_field_0,
  output logic [31:0] o_register_5_bit_field_0,
  output logic [31:0] o_register_6_bit_field_0,
  output logic [31:0] o_register_7_bit_field_0
);

//	altera_conduit_bfm qsys_core_inst_axi4_mst_128_bfm (
//		.sig_araddr  (qsys_core_inst_axi4_mst_128_bfm_conduit_araddr),  // conduit.araddr
//		.sig_arburst (qsys_core_inst_axi4_mst_128_bfm_conduit_arburst), //        .arburst
//		.sig_arlen   (qsys_core_inst_axi4_mst_128_bfm_conduit_arlen),   //        .arlen
//		.sig_arprot  (qsys_core_inst_axi4_mst_128_bfm_conduit_arprot),  //        .arprot
//		.sig_arready (qsys_core_inst_axi4_mst_128_arready),             //        .arready
//		.sig_arsize  (qsys_core_inst_axi4_mst_128_bfm_conduit_arsize),  //        .arsize
//		.sig_arvalid (qsys_core_inst_axi4_mst_128_bfm_conduit_arvalid), //        .arvalid
//		.sig_awaddr  (qsys_core_inst_axi4_mst_128_bfm_conduit_awaddr),  //        .awaddr
//		.sig_awburst (qsys_core_inst_axi4_mst_128_bfm_conduit_awburst), //        .awburst
//		.sig_awlen   (qsys_core_inst_axi4_mst_128_bfm_conduit_awlen),   //        .awlen
//		.sig_awprot  (qsys_core_inst_axi4_mst_128_bfm_conduit_awprot),  //        .awprot
//		.sig_awready (qsys_core_inst_axi4_mst_128_awready),             //        .awready
//		.sig_awsize  (qsys_core_inst_axi4_mst_128_bfm_conduit_awsize),  //        .awsize
//		.sig_awvalid (qsys_core_inst_axi4_mst_128_bfm_conduit_awvalid), //        .awvalid
//		.sig_bready  (qsys_core_inst_axi4_mst_128_bfm_conduit_bready),  //        .bready
//		.sig_bvalid  (qsys_core_inst_axi4_mst_128_bvalid),              //        .bvalid
//		.sig_rdata   (qsys_core_inst_axi4_mst_128_rdata),               //        .rdata
//		.sig_rlast   (qsys_core_inst_axi4_mst_128_rlast),               //        .rlast
//		.sig_rready  (qsys_core_inst_axi4_mst_128_bfm_conduit_rready),  //        .rready
//		.sig_rvalid  (qsys_core_inst_axi4_mst_128_rvalid),              //        .rvalid
//		.sig_wdata   (qsys_core_inst_axi4_mst_128_bfm_conduit_wdata),   //        .wdata
//		.sig_wlast   (qsys_core_inst_axi4_mst_128_bfm_conduit_wlast),   //        .wlast
//		.sig_wready  (qsys_core_inst_axi4_mst_128_wready),              //        .wready
//		.sig_wvalid  (qsys_core_inst_axi4_mst_128_bfm_conduit_wvalid)   //        .wvalid
//	);

	altera_conduit_bfm_0002 qsys_core_inst_axi4_mst_128_reset_bfm (
		.sig_reset (qsys_core_inst_axi4_mst_128_reset_reset)  // conduit.reset
	);

//	altera_conduit_bfm_0003 qsys_core_inst_axi4_mst_16_bfm (
//		.sig_araddr  (qsys_core_inst_axi4_mst_16_bfm_conduit_araddr),  // conduit.araddr
//		.sig_arburst (qsys_core_inst_axi4_mst_16_bfm_conduit_arburst), //        .arburst
//		.sig_arlen   (qsys_core_inst_axi4_mst_16_bfm_conduit_arlen),   //        .arlen
//		.sig_arprot  (qsys_core_inst_axi4_mst_16_bfm_conduit_arprot),  //        .arprot
//		.sig_arready (qsys_core_inst_axi4_mst_16_arready),             //        .arready
//		.sig_arsize  (qsys_core_inst_axi4_mst_16_bfm_conduit_arsize),  //        .arsize
//		.sig_arvalid (qsys_core_inst_axi4_mst_16_bfm_conduit_arvalid), //        .arvalid
//		.sig_awaddr  (qsys_core_inst_axi4_mst_16_bfm_conduit_awaddr),  //        .awaddr
//		.sig_awburst (qsys_core_inst_axi4_mst_16_bfm_conduit_awburst), //        .awburst
//		.sig_awlen   (qsys_core_inst_axi4_mst_16_bfm_conduit_awlen),   //        .awlen
//		.sig_awprot  (qsys_core_inst_axi4_mst_16_bfm_conduit_awprot),  //        .awprot
//		.sig_awready (qsys_core_inst_axi4_mst_16_awready),             //        .awready
//		.sig_awsize  (qsys_core_inst_axi4_mst_16_bfm_conduit_awsize),  //        .awsize
//		.sig_awvalid (qsys_core_inst_axi4_mst_16_bfm_conduit_awvalid), //        .awvalid
//		.sig_bready  (qsys_core_inst_axi4_mst_16_bfm_conduit_bready),  //        .bready
//		.sig_bvalid  (qsys_core_inst_axi4_mst_16_bvalid),              //        .bvalid
//		.sig_rdata   (qsys_core_inst_axi4_mst_16_rdata),               //        .rdata
//		.sig_rlast   (qsys_core_inst_axi4_mst_16_rlast),               //        .rlast
//		.sig_rready  (qsys_core_inst_axi4_mst_16_bfm_conduit_rready),  //        .rready
//		.sig_rvalid  (qsys_core_inst_axi4_mst_16_rvalid),              //        .rvalid
//		.sig_wdata   (qsys_core_inst_axi4_mst_16_bfm_conduit_wdata),   //        .wdata
//		.sig_wlast   (qsys_core_inst_axi4_mst_16_bfm_conduit_wlast),   //        .wlast
//		.sig_wready  (qsys_core_inst_axi4_mst_16_wready),              //        .wready
//		.sig_wvalid  (qsys_core_inst_axi4_mst_16_bfm_conduit_wvalid)   //        .wvalid
//	);

	altera_conduit_bfm_0002 qsys_core_inst_axi4_mst_16_reset_bfm (
		.sig_reset (qsys_core_inst_axi4_mst_16_reset_reset)  // conduit.reset
	);

//	altera_conduit_bfm_0004 qsys_core_inst_axi4lite_slv_0_bfm (
//		.sig_araddr  (qsys_core_inst_axi4lite_slv_0_araddr),              // conduit.araddr
//		.sig_arprot  (qsys_core_inst_axi4lite_slv_0_arprot),              //        .arprot
//		.sig_arready (qsys_core_inst_axi4lite_slv_0_bfm_conduit_arready), //        .arready
//		.sig_arvalid (qsys_core_inst_axi4lite_slv_0_arvalid),             //        .arvalid
//		.sig_awaddr  (qsys_core_inst_axi4lite_slv_0_awaddr),              //        .awaddr
//		.sig_awprot  (qsys_core_inst_axi4lite_slv_0_awprot),              //        .awprot
//		.sig_awready (qsys_core_inst_axi4lite_slv_0_bfm_conduit_awready), //        .awready
//		.sig_awvalid (qsys_core_inst_axi4lite_slv_0_awvalid),             //        .awvalid
//		.sig_bready  (qsys_core_inst_axi4lite_slv_0_bready),              //        .bready
//		.sig_bresp   (qsys_core_inst_axi4lite_slv_0_bfm_conduit_bresp),   //        .bresp
//		.sig_bvalid  (qsys_core_inst_axi4lite_slv_0_bfm_conduit_bvalid),  //        .bvalid
//		.sig_rdata   (qsys_core_inst_axi4lite_slv_0_bfm_conduit_rdata),   //        .rdata
//		.sig_rready  (qsys_core_inst_axi4lite_slv_0_rready),              //        .rready
//		.sig_rresp   (qsys_core_inst_axi4lite_slv_0_bfm_conduit_rresp),   //        .rresp
//		.sig_rvalid  (qsys_core_inst_axi4lite_slv_0_bfm_conduit_rvalid),  //        .rvalid
//		.sig_wdata   (qsys_core_inst_axi4lite_slv_0_wdata),               //        .wdata
//		.sig_wready  (qsys_core_inst_axi4lite_slv_0_bfm_conduit_wready),  //        .wready
//		.sig_wstrb   (qsys_core_inst_axi4lite_slv_0_wstrb),               //        .wstrb
//		.sig_wvalid  (qsys_core_inst_axi4lite_slv_0_wvalid)               //        .wvalid
//	);

	altera_conduit_bfm_0002 qsys_core_inst_axi4lite_slv_0_reset_bfm (
		.sig_reset (qsys_core_inst_axi4lite_slv_0_reset_reset)  // conduit.reset
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (80000000),
		.CLOCK_UNIT (1)
	) qsys_core_inst_clk_bfm (
		.clk (qsys_core_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm_0005 qsys_core_inst_pio_out_bfm (
		.sig_export (qsys_core_inst_pio_out_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) qsys_core_inst_reset_bfm (
		.reset (qsys_core_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (qsys_core_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
